
module conff(
    input wire clock,
    input wire [31:0] bus,
    input wire [31:0] ir,
    input wire con_in,
    output wire con
);

reg con_state;

always @(posedge clock)
begin
    
   
end

endmodule
