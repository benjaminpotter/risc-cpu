module select_encode_logic(input ir, gra, grb, grc, rin, rout, baout, 
                           output [15:0] R_IN, R_OUT
);
	
	
endmodule
									

